
module  FIRST(a,b,c);
input a,b;
output c;
wire d ,clk;
assign c = a+b;

     	 

endmodule